/*
 * datapath.v
 * 
 */
 
/*module datapath(
	input clock,
	input reset,
	input latch_ula,
	input[3:0] ula_operation,
	
	inout[7:0] data_bus
);

wire[7:0]  register_operand;
wire[15:0] ula_result;

ula m_ula(clock, reset, register_operand, data_bus, ula_operation, ula_result);

endmodule
*/
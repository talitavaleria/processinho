/*
 * program_counter.v
 * 
 */

module program_counter(
	input clock
)




endmodule
